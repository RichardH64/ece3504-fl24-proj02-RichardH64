////////////////////////////////////////////////////////////////
//  Filename     : mips.v
//  Module       : MIPS
//  Author       : L. Nazhand-Ali
//  Modified by  : C. Patterson, R. Harrison (18 Nov 2024)
//  Description  : single cycle MIPS 
//   
//     The top module of the single cycle MIPS is presented in this
//  file. You need to edit this module to complete the data path for
//  some of the instructions in your project.


module MIPS(clk, reset);

   input clk;
   input reset;

   // instruction and PC related wires
   wire [31:0] instruction;
   wire [31:0] PCplus4;
   wire [31:0]    //===Added Modules (18 Nov 2024)===//
   // instantiation of a 32-bit 2-bit left shifter used for shifting the branch offset for branch target address calculation
   SHIFT2 shift2
      (
      .word_out(immShifted),
      .word_in(immExtended)
      );
      
   // instantiation of a 32-bit adder used for computing branch target
   ADDER32 branchAdder
     (
      .result_out(branchPC),
      .a_in(PCplus4), 
      .b_in(immShifted)
      );
   
   // instantiation of a 32-bit MUX used for selecting between PC+4 and branch address as the nextPC
   MUX32_2X1 branchMux
     (
      .value_out(nextPC),
      .value0_in(PCplus4), 
      .value1_in(branchPC), 
      .select_in(jump | branch)
      );;
   
   // decoder related wires
   wire [5:0]  op, func;
   wire [4:0]  rs, rt, rd, shft;
   wire [15:0] imm16;
   wire [25:0] target;
   
   // control related wires
   wire        regWrite, regDst;
   wire        memRead, memWrite, memToReg;
   wire        extCntrl, ALUSrc;
   wire [3:0]  ALUCntrl;
   wire        branch, jump;

   // ALU related wires
   wire [31:0] A, B, ALUout;
   wire        zero;

   // register file related wires
   wire [31:0] regData2;
   wire [4:0]  regDstAddr;

   // immediate related wires
   wire [31:0] immExtended;

   ///////////////////////////////////////////////
   // Put your new wires below this line
   wire [31:0] immShifted;
   wire [31:0] targetShifted;
   wire [31:0] branchAddr;
   wire [31:0] jumpAddr;
   wire [31:0] branchJump
   wire [31:0] nextPC;
   wire [31:0] finalPC;
   
   //////////////////////////////////////////////
   

   // instantiation of instruction memory
   IMEM	imem
     (
      .instruction_out(instruction),
      .address_in(PC)
      );


   // instantiation of register file
   REG_FILE reg_file
     (
      .clk(clk),
      .data1_out(A),
      .data2_out(regData2),
      .readAddr1_in(rs),
      .readAddr2_in(rt),
      .writeAddr_in(regDstAddr),
      .writeData_in(ALUout),
      .writeCntrl_in(regWrite)
      );

   // instantiation of PC register //===Modified (18 Nov 2024)===//
   PC_REG pc_reg
     (
      .clk(clk),
      .reset(reset),
      .PC_out(PC),
      .PC_in(finalPC)
      );

   // instantiation of the decoder
   MIPS_DECODE	mips_decode
     (
      .instruction_in(instruction), 
      .op_out(op), 
      .func_out(func), 
      .rs_out(rs), 
      .rt_out(rt), 
      .rd_out(rd), 
      .shft_out(shft), 
      .imm16_out(imm16), 
      .target_out(target)
      );

   // instantiation of the control unit
   MIPS_CONTROL mips_control
     (
      .op_in(op),
      .func_in(func),
      .branch_out(branch), 
      .regWrite_out(regWrite), 
      .regDst_out(regDst), 
      .extCntrl_out(extCntrl), 
      .ALUSrc_out(ALUSrc), 
      .ALUCntrl_out(ALUCntrl), 
      .memWrite_out(memWrite),
      .memRead_out(memRead),
      .memToReg_out(memToReg), 
      .jump_out(jump)
      );

   // instantiation of the ALU
   MIPS_ALU mips_alu
     (
      .ALUCntrl_in(ALUCntrl), 
      .A_in(A), 
      .B_in(B), 
      .ALU_out(ALUout), 
      .zero_out(zero)
      );

   // instantiation of the sign/zero extender
   EXTEND extend
     (
      .word_out(immExtended),
      .halfWord_in(imm16),
      .extendCntrl_in(extCntrl)
      );

   // instantiation of a 32-bit adder used for computing PC+4
   ADDER32 plus4Adder
     (
      .result_out(PCplus4),
      .a_in(32'd4), 
      .b_in(PC)
      );

   // instantiation of a 32-bit MUX used for selecting between immediate and register as the second source of ALU
   MUX32_2X1 aluMux
     (
      .value_out(B),
      .value0_in(regData2), 
      .value1_in(immExtended), 
      .select_in(ALUSrc)
      );

   // instantiation of a 5-bit MUX used for selecting between RT or RD as the destination address of the operation
   MUX5_2X1 regMUX 
     (
      .value_out(regDstAddr),
      .value0_in(rt),
      .value1_in(rd),
      .select_in(regDst)
      );
   
   //===Added Modules (18 Nov 2024)===//
   // instantiation of a 32-bit 2-bit shift left used for shifting the target for jump target address calculation
   SHIFT2 jumpShift (
       .word_out(targetShifted),
       .word_in({6'b0, target_out})
   );

   // Concatenate upper 4 bits of PC+4 with shifted target
   assign jumpAddr = {PCplus4[31:28], targetShifted[27:0]};
   
   // instantiation of a 32-bit 2-bit shift left used for shifting the branch offset for branch target address calculation
   SHIFT2 immShift
      (
      .word_out(immShifted),
      .word_in(immExtended)
      );
   
   // instantiation of a 32-bit adder used for computing branch target
   ADDER32 branchAdder
     (
      .result_out(branchPC),
      .a_in(PCplus4), 
      .b_in(immShifted)
      );
   
   // instantiation of a 32-bit MUX used for selecting between PC+4 and branch address as the nextPC
   MUX32_2X1 branchMux
     (
      .value_out(nextPC),
      .value0_in(PCplus4), 
      .value1_in(branchPC), 
      .select_in(branch)
      );
   
   // instantiation of a 32-bit MUX used for selecting between nextPC (PC+4 or branchAddr) and jumAddr as the finalPC
   MUX32_2X1 jumpMux
     (
      .value_out(finalPC),
      .value0_in(nextPC), 
      .value1_in(jumpAddr), 
      .select_in(jump)
      );
endmodule
